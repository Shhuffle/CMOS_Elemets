** sch_path: /home/safal/projects/CMOS_Elemets/Schematic/VoltageDivider.sch
**.subckt VoltageDivider
XR1 V_Out V_In Gnd sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR2 net1 V_Out Gnd sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR3 net2 net1 Gnd sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR4 net3 net2 Gnd sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR5 Gnd net3 Gnd sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR6 net4 net5 Gnd sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
XR7 net6 net7 Gnd sky130_fd_pr__res_xhigh_po_0p35 L=0.35 mult=1 m=1
**.ends
.GLOBAL Gnd
.end
