magic
tech sky130A
timestamp 1748943440
<< psubdiff >>
rect 28261 13449 28361 13451
rect 28015 13377 28361 13449
rect 28015 13294 28080 13377
rect 28198 13294 28361 13377
rect 28015 13238 28361 13294
<< psubdiffcont >>
rect 28080 13294 28198 13377
<< xpolycontact >>
rect 26629 13885 26664 14105
rect 26629 13319 26664 13539
rect 26709 13885 26744 14105
rect 26709 13319 26744 13539
rect 26799 13884 26834 14104
rect 26799 13318 26834 13538
rect 26887 13886 26922 14106
rect 26887 13320 26922 13540
rect 26977 13885 27012 14105
rect 26977 13319 27012 13539
rect 27053 13886 27088 14106
rect 27053 13320 27088 13540
rect 27143 13885 27178 14105
rect 27143 13319 27178 13539
<< xpolyres >>
rect 26629 13539 26664 13885
rect 26709 13539 26744 13885
rect 26799 13538 26834 13884
rect 26887 13540 26922 13886
rect 26977 13539 27012 13885
rect 27053 13540 27088 13886
rect 27143 13539 27178 13885
<< locali >>
rect 26525 14046 26567 14063
rect 26594 14046 26629 14062
rect 26599 13943 26629 14046
rect 26594 13924 26629 13943
rect 26664 13924 26665 14062
rect 26834 13886 26887 14104
rect 27012 13886 27053 14104
rect 26744 13538 26804 13539
rect 26744 13321 26799 13538
rect 26922 13320 26977 13537
rect 26919 13319 26977 13320
rect 27049 13320 27053 13411
rect 27088 13320 27091 13411
rect 27049 13235 27091 13320
rect 28040 13378 28229 13405
rect 28040 13294 28079 13378
rect 28199 13294 28229 13378
rect 28040 13269 28229 13294
<< viali >>
rect 26494 13943 26599 14046
rect 28079 13377 28199 13378
rect 28079 13294 28080 13377
rect 28080 13294 28198 13377
rect 28198 13294 28199 13377
rect 27018 13132 27123 13235
<< metal1 >>
rect 26489 14046 26606 14052
rect 26489 13943 26494 14046
rect 26599 13943 26606 14046
rect 26489 13937 26606 13943
rect 27961 13388 28327 13405
rect 27961 13278 28066 13388
rect 28213 13278 28327 13388
rect 27961 13269 28327 13278
rect 28042 13267 28228 13269
rect 27013 13235 27130 13241
rect 27013 13132 27018 13235
rect 27123 13132 27130 13235
rect 27013 13126 27130 13132
<< via1 >>
rect 26500 13951 26590 14039
rect 28066 13378 28213 13388
rect 28066 13294 28079 13378
rect 28079 13294 28199 13378
rect 28199 13294 28213 13378
rect 28066 13278 28213 13294
rect 27024 13140 27114 13228
<< metal2 >>
rect 26497 14039 26594 14042
rect 26497 13951 26500 14039
rect 26590 13951 26594 14039
rect 26497 13947 26594 13951
rect 28055 13388 28223 13399
rect 28055 13278 28066 13388
rect 28213 13278 28223 13388
rect 27021 13228 27118 13231
rect 27021 13140 27024 13228
rect 27114 13140 27118 13228
rect 28055 13227 28090 13278
rect 28199 13227 28223 13278
rect 28055 13173 28223 13227
rect 27021 13136 27118 13140
<< via2 >>
rect 26503 13954 26587 14036
rect 28090 13278 28199 13345
rect 27027 13143 27111 13225
rect 28090 13227 28199 13278
<< metal3 >>
rect 26480 14036 26615 14042
rect 26480 13954 26503 14036
rect 26587 13954 26615 14036
rect 26480 13951 26615 13954
rect 26485 13949 26607 13951
rect 27195 13505 28300 14598
rect 27981 13451 28300 13505
rect 27981 13345 28322 13451
rect 27004 13225 27139 13231
rect 27004 13143 27027 13225
rect 27111 13143 27139 13225
rect 27981 13227 28090 13345
rect 28199 13238 28322 13345
rect 28199 13227 28300 13238
rect 27981 13219 28300 13227
rect 27004 13140 27139 13143
rect 27009 13138 27131 13140
rect 28082 13020 28216 13219
<< via3 >>
rect 26508 13957 26582 14030
rect 27032 13146 27106 13219
<< mimcap >>
rect 27295 14002 28186 14498
rect 27295 13700 27394 14002
rect 27633 13700 28186 14002
rect 27295 13607 28186 13700
<< mimcapcontact >>
rect 27394 13700 27633 14002
<< metal4 >>
rect 26477 14052 26623 14061
rect 26413 14030 26623 14052
rect 26413 13957 26508 14030
rect 26582 13957 26623 14030
rect 26413 13937 26623 13957
rect 26477 13925 26623 13937
rect 27375 14002 27652 14029
rect 27375 13700 27394 14002
rect 27633 13700 27652 14002
rect 27375 13250 27652 13700
rect 26970 13222 27652 13250
rect 26970 13219 27649 13222
rect 26970 13146 27032 13219
rect 27106 13146 27649 13219
rect 26970 13096 27649 13146
rect 26970 13094 27407 13096
<< labels >>
rlabel metal4 27496 13238 27496 13238 1 V_Out
port 1 n
rlabel metal4 26414 13991 26414 13991 3 V_In
port 2 e
rlabel psubdiff 28359 13328 28359 13328 7 Gnd
<< end >>
