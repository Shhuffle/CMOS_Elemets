* SPICE3 file created from NMOS.ext - technology: sky130A

X0 a_10_0# a_n20_n26# a_n74_0# a_n186_n2# sky130_fd_pr__nfet_01v8 ad=0.1215 pd=1.44 as=0.1215 ps=1.44 w=0.45 l=0.15
